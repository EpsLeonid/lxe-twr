library ieee;
use ieee.std_logic_1164.all;

package constants is
	
	constant DATA_WIDTH : integer := 12;
	constant DATA_WIDTH_DIV_2 : integer := DATA_WIDTH/2;
	
end constants;

package body constants is
end constants;

